module coprocessor (input logic clk, Start,
                    input logic [31:0] WriteData,
                    output logic done,
                    output logic [31:0] ReadData);

// stuff here


endmodule
