module coprocessor (input logic clk, Start,
                    input logic [31:0] WDFinal,
                    output logic copDone,
                    output logic [31:0] AnsData);

// stuff here


endmodule